module hsync(
    clk,
    reset,
    hPixel,
    display_active,
    hsync
);

input clk, reset;
output [6:0] hPixel;
output display_active;
output hsync;

reg [6:0] hPixel;
reg rgb_active;
reg display_active;
reg hsync;


reg [2:0] currentState, nextState;

reg [12:0] state_counter;
reg reset_state_counter;

reg [5:0] pixel_counter;
reg pixel_enable;

parameter OFF=3'b000,
          HSYNC_PULSE_WIDTH=3'b001,
          BACK_PORCH=3'b010,
          DISPLAY=3'b011,
          FRONT_PORCH=3'b100;

parameter PULSE_WIDTH_TIME=384,
          BACK_PORCH_TIME=192,
          DISPLAY_TIME=2560,
          FRONT_PORCH_TIME=64;

/*an always to handle the state_counter.
The counter gets to 0 when reset is asserted
or when the hsync gets to the PULSE_WIDTH
state again where the reset_state_counter
reset the counter*/
always@(posedge clk or posedge reset)
    begin
        if(reset) begin
            state_counter<=13'b0;
        end
        else if(reset_state_counter)
            state_counter<=13'b0;
        else
        state_counter<=state_counter+1;
    end

always@(posedge clk or posedge reset)
    begin
        if(reset)
            pixel_counter<=4'b0000;
         else begin
            
         
        if(pixel_enable) begin
            pixel_counter<=pixel_counter+1;
            if(pixel_counter==19) begin
                hPixel<=hPixel+1;
                pixel_counter<=4'b0000;
            end
        end
        else begin
            pixel_counter<=4'b0000;
            hPixel<=1'b0;
        end
        end

    end

/*always that changes the states*/
always@(posedge clk or posedge reset)
    begin
        if(reset)
            currentState<=OFF;
        else
            currentState<=nextState;
    end

always@(currentState or state_counter)
    begin
        nextState=currentState;
        hsync=1'b0;
        display_active=1'b0;
        reset_state_counter=1'b0;
        pixel_enable=1'b0;

        case(currentState)
            OFF: begin
                hsync=1'b0;
                display_active=1'b0;
                reset_state_counter=1'b1;
                pixel_enable=1'b0;
                
                nextState=HSYNC_PULSE_WIDTH;
            end

            HSYNC_PULSE_WIDTH: begin
                hsync=1'b0;
                display_active=1'b0;
                reset_state_counter=1'b0;
                pixel_enable=1'b0;

                if(state_counter==PULSE_WIDTH_TIME-1) begin //count to 3.84us (92 cycles)
                    nextState=BACK_PORCH;
                    // reset_state_counter=1'b0;
                end
                else begin
                    nextState=HSYNC_PULSE_WIDTH;
                    // reset_state_counter=1'b0;
                end
            end

            BACK_PORCH: begin
                hsync=1'b1;
                display_active=1'b0;
                reset_state_counter=1'b0;
                pixel_enable=1'b0;

                if(state_counter==(PULSE_WIDTH_TIME+BACK_PORCH)-1)//count 3.84us+1.92us (192+96 cycles)
                    nextState=DISPLAY;
                else
                    nextState=BACK_PORCH;
            end

            DISPLAY: begin
                hsync=1'b1;
                display_active=1'b1;
                reset_state_counter=1'b0;
                pixel_enable=1'b1;

                if(state_counter==(PULSE_WIDTH_TIME+BACK_PORCH+DISPLAY_TIME)-1)//count 3.84us+1.92us+25.6us(192+96+1280 cycles)
                    nextState=FRONT_PORCH;
                else
                    nextState=DISPLAY;
            end

            FRONT_PORCH: begin
                hsync=1'b1;
                display_active=1'b0;
                reset_state_counter=1'b0;
                pixel_enable=1'b0;

                if(state_counter==(PULSE_WIDTH_TIME+BACK_PORCH+DISPLAY_TIME+FRONT_PORCH_TIME)-1) begin//count 3.84us+1.92us+25.6us+0.64us(192+96+1280+32 cycles)
                    nextState=HSYNC_PULSE_WIDTH;
                    reset_state_counter=1'b1;
                end
                else
                    nextState=FRONT_PORCH;
            end
        endcase
    end
endmodule