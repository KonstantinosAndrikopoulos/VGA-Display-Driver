//  RAMB18E1   : In order to incorporate this function into the design,
//   Verilog   : the following instance declaration needs to be placed
//  instance   : in the body of the design code.  The instance name
// declaration : (RAMB18E1_inst) and/or the port declarations within the
//    code     : parenthesis may be changed to properly reference and
//             : connect this function to the design.  All inputs
//             : and outputs must be connected.

//  <-----Cut code below this line---->

   // RAMB18E1: 18K-bit Configurable Synchronous Block RAM
   //           Artix-7
   // Xilinx HDL Language Template, version 2018.3

    module VRAM (
        clk,
        reset,
        read_address,
        read_enable,
        rgb,
        write_enable,
        R_write_data_low,
        R_write_data_upper,
        G_write_data_low,
        G_write_data_upper,
        B_write_data_low,
        B_write_data_upper,
        write_address
    );

    input reset, clk;
    
    //128x96 VRAM that means we need 2^7 and also 2^7 so {}
    input [13:0] read_address;
    input read_enable;
    
    //rgb[2]=red, rgb[1]=green, rgb[0]=blue
    output [2:0] rgb;

    //write inputs
    input [3:0] write_enable;
    input [13:0] write_address;

    input [15:0]  R_write_data_low, R_write_data_upper, G_write_data_low, G_write_data_upper, B_write_data_low, B_write_data_upper;

    wire [15:0] doa_data_red, doa_data_green, doa_data_blue;

   assign rgb[2] = doa_data_red[0]; // Assuming you need the LSB
   assign rgb[1] = doa_data_green[0];
   assign rgb[0] = doa_data_blue[0];

   RAMB18E1 #(
      // Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE" 
      .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
      // Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
      .SIM_COLLISION_CHECK("ALL"),
      // DOA_REG, DOB_REG: Optional output register (0 or 1)
      .DOA_REG(0),
      .DOB_REG(0),
      // INITP_00 to INITP_07: Initial contents of parity memory array
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // INIT_00 to INIT_3F: Initial contents of data memory array
      .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),


      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF), 
      .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_24(256'hFFFFFFFFF000000FFFFFF000000FFFFF_FFFFFFFFF000000FFFFFF000000FFFFF),
      .INIT_25(256'hFFFFFFFFF000000FFFFFF000000FFFFF_FFFFFFFFF000000FFFFFF000000FFFFF),
      .INIT_26(256'hFFFFFFFFF000000FFFFFF000000FFFFF_FFFFFFFFF000000FFFFFF000000FFFFF),
      .INIT_27(256'hFFFFFFFFF000000FFFFFF000000FFFFF_FFFFFFFFF000000FFFFFF000000FFFFF),
      .INIT_28(256'h000000FFF000000FFFFFF00000000000_000000FFF000000FFFFFF00000000000),
      .INIT_29(256'h000000FFF000000FFFFFF00000000000_000000FFF000000FFFFFF00000000000),
      .INIT_2A(256'h000000FFF000000FFFFFF00000000000_000000FFF000000FFFFFF00000000000),
      .INIT_2B(256'h000000FFF000000FFFFFF00000000000_000000FFF000000FFFFFF00000000000),
      .INIT_2C(256'hFFFFFFFFF000000FFFFFF000000FFFFF_FFFFFFFFF000000FFFFFF000000FFFFF),
      .INIT_2D(256'hFFFFFFFFF000000FFFFFF000000FFFFF_FFFFFFFFF000000FFFFFF000000FFFFF),
      .INIT_2E(256'hFFFFFFFFF000000FFFFFF000000FFFFF_FFFFFFFFF000000FFFFFF000000FFFFF),
      .INIT_2F(256'hFFFFFFFFF000000FFFFFF000000FFFFF_FFFFFFFFF000000FFFFFF000000FFFFF),
      .INIT_30(256'h00000FFFFF000000000000000FFFFF000000000000000FFFFF00000000000000),
      .INIT_31(256'h00000FFFFF000000000000000FFFFF000000000000000FFFFF00000000000000),
      .INIT_32(256'h00000FFFFF000000000000000FFFFF000000000000000FFFFF00000000000000),
      .INIT_33(256'h00000FFFFF000000000000000FFFFF000000000000000FFFFF00000000000000),
      .INIT_34(256'hFFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFF),
      .INIT_35(256'hFFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFF),
      .INIT_36(256'hFFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFF),
      .INIT_37(256'hFFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFF),
      .INIT_38(256'h00000FFFFF000000000000000FFFFF000000000000000FFFFF00000000000000),
      .INIT_39(256'h00000FFFFF000000000000000FFFFF000000000000000FFFFF00000000000000),
      .INIT_3A(256'h00000FFFFF000000000000000FFFFF000000000000000FFFFF00000000000000),
      .INIT_3B(256'h00000FFFFF000000000000000FFFFF000000000000000FFFFF00000000000000),
      .INIT_3C(256'hFFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFF),
      .INIT_3D(256'hFFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFF),
      .INIT_3E(256'hFFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFF),
      .INIT_3F(256'hFFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFF),
      // INIT_A, INIT_B: Initial values on output ports
      .INIT_A(18'h00000),
      .INIT_B(18'h00000),
      // Initialization File: RAM initialization file
      .INIT_FILE("NONE"),
      // RAM Mode: "SDP" or "TDP" 
      .RAM_MODE("SDP"),
      // READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
      .READ_WIDTH_A(1),                                                                 // 0-72
      .READ_WIDTH_B(0),                                                                 // 0-18
      .WRITE_WIDTH_A(0),                                                                // 0-18
      .WRITE_WIDTH_B(36),                                                                // 0-72
      // RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
      .RSTREG_PRIORITY_A("RSTREG"),
      .RSTREG_PRIORITY_B("RSTREG"),
      // SRVAL_A, SRVAL_B: Set/reset value for output
      .SRVAL_A(18'h00000),
      .SRVAL_B(18'h00000),
      // Simulation Device: Must be set to "7SERIES" for simulation behavior
      .SIM_DEVICE("7SERIES"),
      // WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
      .WRITE_MODE_A("WRITE_FIRST"),
      .WRITE_MODE_B("WRITE_FIRST")
   )
   VRAM_RED (
      // Port A Data: 16-bit (each) output: Port A data
      .DOADO(doa_data_red),                 // 16-bit output: A port data/LSB data
      .DOPADOP(),             // 2-bit output: A port parity/LSB parity
      // Port B Data: 16-bit (each) output: Port B data
      .DOBDO(),                 // 16-bit output: B port data/MSB data
      .DOPBDOP(),             // 2-bit output: B port parity/MSB parity
      // Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals (read port
      // when RAM_MODE="SDP")
      .ADDRARDADDR(read_address),     // 14-bit input: A port address/Read address
      .CLKARDCLK(clk),         // 1-bit input: A port clock/Read clock
      .ENARDEN(read_enable),             // 1-bit input: A port enable/Read enable
      .REGCEAREGCE(1'b0),     // 1-bit input: A port register enable/Register enable
      .RSTRAMARSTRAM(reset), // 1-bit input: A port set/reset
      .RSTREGARSTREG(1'b0), // 1-bit input: A port register set/reset
      .WEA(),                     // 2-bit input: A port write enable
      // Port A Data: 16-bit (each) input: Port A data
      .DIADI(R_write_data_low),                 // 16-bit input: A port data/LSB data
      .DIPADIP(),             // 2-bit input: A port parity/LSB parity
      // Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals (write port
      // when RAM_MODE="SDP")
      .ADDRBWRADDR(write_address),     // 14-bit input: B port address/Write address
      .CLKBWRCLK(clk),         // 1-bit input: B port clock/Write clock
      .ENBWREN(1'b1),             // 1-bit input: B port enable/Write enable
      .REGCEB(),               // 1-bit input: B port register enable
      .RSTRAMB(),             // 1-bit input: B port set/reset
      .RSTREGB(),             // 1-bit input: B port register set/reset
      .WEBWE(write_enable),                 // 4-bit input: B port write enable/Write enable
      // Port B Data: 16-bit (each) input: Port B data
      .DIBDI(R_write_data_upper),                 // 16-bit input: B port data/MSB data
      .DIPBDIP()              // 2-bit input: B port parity/MSB parity
   );

    RAMB18E1 #(
      // Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE" 
      .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
      // Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
      .SIM_COLLISION_CHECK("ALL"),
      // DOA_REG, DOB_REG: Optional output register (0 or 1)
      .DOA_REG(0),
      .DOB_REG(0),
      // INITP_00 to INITP_07: Initial contents of parity memory array
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // INIT_00 to INIT_3F: Initial contents of data memory array
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),


      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_24(256'hFFFFFF000FFF000FFF000FFF000FFFFF_FFFFFF000FFF000FFF000FFF000FFFFF),
      .INIT_25(256'hFFFFFF000FFF000FFF000FFF000FFFFF_FFFFFF000FFF000FFF000FFF000FFFFF),
      .INIT_26(256'hFFFFFF000FFF000FFF000FFF000FFFFF_FFFFFF000FFF000FFF000FFF000FFFFF),
      .INIT_27(256'hFFFFFF000FFF000FFF000FFF000FFFFF_FFFFFF000FFF000FFF000FFF000FFFFF),
      .INIT_28(256'h000000000FFF000FFF000FFF00000000_000000000FFF000FFF000FFF00000000),
      .INIT_29(256'h000000000FFF000FFF000FFF00000000_000000000FFF000FFF000FFF00000000),
      .INIT_2A(256'h000000000FFF000FFF000FFF00000000_000000000FFF000FFF000FFF00000000),
      .INIT_2B(256'h000000000FFF000FFF000FFF00000000_000000000FFF000FFF000FFF00000000),
      .INIT_2C(256'hFFFFFF000FFF000FFF000FFF000FFFFF_FFFFFF000FFF000FFF000FFF000FFFFF),
      .INIT_2D(256'hFFFFFF000FFF000FFF000FFF000FFFFF_FFFFFF000FFF000FFF000FFF000FFFFF),
      .INIT_2E(256'hFFFFFF000FFF000FFF000FFF000FFFFF_FFFFFF000FFF000FFF000FFF000FFFFF),
      .INIT_2F(256'hFFFFFF000FFF000FFF000FFF000FFFFF_FFFFFF000FFF000FFF000FFF000FFFFF),
      .INIT_30(256'h0000000000FFFFF000000000000000FFFFF000000000000000FFFFF000000000),
      .INIT_31(256'h0000000000FFFFF000000000000000FFFFF000000000000000FFFFF000000000),
      .INIT_32(256'h0000000000FFFFF000000000000000FFFFF000000000000000FFFFF000000000),
      .INIT_33(256'h0000000000FFFFF000000000000000FFFFF000000000000000FFFFF000000000),
      .INIT_34(256'hFFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFF),
      .INIT_35(256'hFFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFF),
      .INIT_36(256'hFFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFF),
      .INIT_37(256'hFFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFF),
      .INIT_38(256'h0000000000FFFFF000000000000000FFFFF000000000000000FFFFF000000000),
      .INIT_39(256'h0000000000FFFFF000000000000000FFFFF000000000000000FFFFF000000000),
      .INIT_3A(256'h0000000000FFFFF000000000000000FFFFF000000000000000FFFFF000000000),
      .INIT_3B(256'h0000000000FFFFF000000000000000FFFFF000000000000000FFFFF000000000),
      .INIT_3C(256'hFFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFF),
      .INIT_3D(256'hFFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFF),
      .INIT_3E(256'hFFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFF),
      .INIT_3F(256'hFFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFFF00000FFFF),
      // INIT_A, INIT_B: Initial values on output ports
      .INIT_A(1'b0),
      .INIT_B(18'h00000),
      // Initialization File: RAM initialization file
      .INIT_FILE("NONE"),
      // RAM Mode: "SDP" or "TDP" 
      .RAM_MODE("SDP"),
      // READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
      .READ_WIDTH_A(1),                                                                 // 0-72
      .READ_WIDTH_B(0),                                                                 // 0-18
      .WRITE_WIDTH_A(0),                                                                // 0-18
      .WRITE_WIDTH_B(36),                                                                // 0-72
      // RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
      .RSTREG_PRIORITY_A("RSTREG"),
      .RSTREG_PRIORITY_B("RSTREG"),
      // SRVAL_A, SRVAL_B: Set/reset value for output
      .SRVAL_A(18'h00000),
      .SRVAL_B(18'h00000),
      // Simulation Device: Must be set to "7SERIES" for simulation behavior
      .SIM_DEVICE("7SERIES"),
      // WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
      .WRITE_MODE_A("WRITE_FIRST"),
      .WRITE_MODE_B("WRITE_FIRST")
   )
   VRAM_GREEN (
      // Port A Data: 16-bit (each) output: Port A data
      .DOADO(doa_data_green),                 // 16-bit output: A port data/LSB data
      .DOPADOP(),             // 2-bit output: A port parity/LSB parity
      // Port B Data: 16-bit (each) output: Port B data
      .DOBDO(),                 // 16-bit output: B port data/MSB data
      .DOPBDOP(),             // 2-bit output: B port parity/MSB parity
      // Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals (read port
      // when RAM_MODE="SDP")
      .ADDRARDADDR(read_address),     // 14-bit input: A port address/Read address
      .CLKARDCLK(clk),         // 1-bit input: A port clock/Read clock
      .ENARDEN(read_enable),             // 1-bit input: A port enable/Read enable
      .REGCEAREGCE(1'b0),     // 1-bit input: A port register enable/Register enable
      .RSTRAMARSTRAM(reset), // 1-bit input: A port set/reset
      .RSTREGARSTREG(1'b0), // 1-bit input: A port register set/reset
      .WEA(),                     // 2-bit input: A port write enable
      // Port A Data: 16-bit (each) input: Port A data
      .DIADI(G_write_data_low),                 // 16-bit input: A port data/LSB data
      .DIPADIP(),             // 2-bit input: A port parity/LSB parity
      // Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals (write port
      // when RAM_MODE="SDP")
      .ADDRBWRADDR(write_address),     // 14-bit input: B port address/Write address
      .CLKBWRCLK(clk),         // 1-bit input: B port clock/Write clock
      .ENBWREN(1'b1),             // 1-bit input: B port enable/Write enable
      .REGCEB(),               // 1-bit input: B port register enable
      .RSTRAMB(),             // 1-bit input: B port set/reset
      .RSTREGB(),             // 1-bit input: B port register set/reset
      .WEBWE(write_enable),                 // 4-bit input: B port write enable/Write enable
      // Port B Data: 16-bit (each) input: Port B data
      .DIBDI(G_write_data_upper),                 // 16-bit input: B port data/MSB data
      .DIPBDIP()              // 2-bit input: B port parity/MSB parity
   );

       RAMB18E1 #(
      // Address Collision Mode: "PERFORMANCE" or "DELAYED_WRITE" 
      .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
      // Collision check: Values ("ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE")
      .SIM_COLLISION_CHECK("ALL"),
      // DOA_REG, DOB_REG: Optional output register (0 or 1)
      .DOA_REG(0),
      .DOB_REG(0),
      // INITP_00 to INITP_07: Initial contents of parity memory array
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // INIT_00 to INIT_3F: Initial contents of data memory array
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),


      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_24(256'hFFFFFF000000FFFFFF000000FFFFFFFF_FFFFFF000000FFFFFF000000FFFFFFFF),
      .INIT_25(256'hFFFFFF000000FFFFFF000000FFFFFFFF_FFFFFF000000FFFFFF000000FFFFFFFF),
      .INIT_26(256'hFFFFFF000000FFFFFF000000FFFFFFFF_FFFFFF000000FFFFFF000000FFFFFFFF),
      .INIT_27(256'hFFFFFF000000FFFFFF000000FFFFFFFF_FFFFFF000000FFFFFF000000FFFFFFFF),
      .INIT_28(256'h000000000000FFFFFF000000FFF00000_000000000000FFFFFF000000FFF00000),
      .INIT_29(256'h000000000000FFFFFF000000FFF00000_000000000000FFFFFF000000FFF00000),
      .INIT_2A(256'h000000000000FFFFFF000000FFF00000_000000000000FFFFFF000000FFF00000),
      .INIT_2B(256'h000000000000FFFFFF000000FFF00000_000000000000FFFFFF000000FFF00000),
      .INIT_2C(256'hFFFFFF000000FFFFFF000000FFFFFFFF_FFFFFF000000FFFFFF000000FFFFFFFF),
      .INIT_2D(256'hFFFFFF000000FFFFFF000000FFFFFFFF_FFFFFF000000FFFFFF000000FFFFFFFF),
      .INIT_2E(256'hFFFFFF000000FFFFFF000000FFFFFFFF_FFFFFF000000FFFFFF000000FFFFFFFF),
      .INIT_2F(256'hFFFFFF000000FFFFFF000000FFFFFFFF_FFFFFF000000FFFFFF000000FFFFFFFF),
      .INIT_30(256'h000000000000000FFFFF000000000000000FFFFF000000000000000FFFFF0000),
      .INIT_31(256'h000000000000000FFFFF000000000000000FFFFF000000000000000FFFFF0000),
      .INIT_32(256'h000000000000000FFFFF000000000000000FFFFF000000000000000FFFFF0000),
      .INIT_33(256'h000000000000000FFFFF000000000000000FFFFF000000000000000FFFFF0000),
      .INIT_34(256'hFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFF),
      .INIT_35(256'hFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFF),
      .INIT_36(256'hFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFF),
      .INIT_37(256'hFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFF),
      .INIT_38(256'h000000000000000FFFFF000000000000000FFFFF000000000000000FFFFF0000),
      .INIT_39(256'h000000000000000FFFFF000000000000000FFFFF000000000000000FFFFF0000),
      .INIT_3A(256'h000000000000000FFFFF000000000000000FFFFF000000000000000FFFFF0000),
      .INIT_3B(256'h000000000000000FFFFF000000000000000FFFFF000000000000000FFFFF0000),
      .INIT_3C(256'hFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFF),
      .INIT_3D(256'hFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFF),
      .INIT_3E(256'hFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFF),
      .INIT_3F(256'hFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFFF0000000000FFFFFFFFF),
      // INIT_A, INIT_B: Initial values on output ports
      .INIT_A(18'h00000),
      .INIT_B(18'h00000),
      // Initialization File: RAM initialization file
      .INIT_FILE("NONE"),
      // RAM Mode: "SDP" or "TDP" 
      .RAM_MODE("SDP"),
      // READ_WIDTH_A/B, WRITE_WIDTH_A/B: Read/write width per port
      .READ_WIDTH_A(1),                                                                 // 0-72
      .READ_WIDTH_B(0),                                                                 // 0-18
      .WRITE_WIDTH_A(0),                                                                // 0-18
      .WRITE_WIDTH_B(36),                                                                // 0-72
      // RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
      .RSTREG_PRIORITY_A("RSTREG"),
      .RSTREG_PRIORITY_B("RSTREG"),
      // SRVAL_A, SRVAL_B: Set/reset value for output
      .SRVAL_A(18'h00000),
      .SRVAL_B(18'h00000),
      // Simulation Device: Must be set to "7SERIES" for simulation behavior
      .SIM_DEVICE("7SERIES"),
      // WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
      .WRITE_MODE_A("WRITE_FIRST"),
      .WRITE_MODE_B("WRITE_FIRST")
   )
   VRAM_BLUE (
      // Port A Data: 16-bit (each) output: Port A data
      .DOADO(doa_data_blue),                 // 16-bit output: A port data/LSB data
      .DOPADOP(),             // 2-bit output: A port parity/LSB parity
      // Port B Data: 16-bit (each) output: Port B data
      .DOBDO(),                 // 16-bit output: B port data/MSB data
      .DOPBDOP(),             // 2-bit output: B port parity/MSB parity
      // Port A Address/Control Signals: 14-bit (each) input: Port A address and control signals (read port
      // when RAM_MODE="SDP")
      .ADDRARDADDR(read_address),     // 14-bit input: A port address/Read address
      .CLKARDCLK(clk),         // 1-bit input: A port clock/Read clock
      .ENARDEN(read_enable),             // 1-bit input: A port enable/Read enable
      .REGCEAREGCE(1'b0),     // 1-bit input: A port register enable/Register enable
      .RSTRAMARSTRAM(reset), // 1-bit input: A port set/reset
      .RSTREGARSTREG(1'b0), // 1-bit input: A port register set/reset
      .WEA(),                     // 2-bit input: A port write enable
      // Port A Data: 16-bit (each) input: Port A data
      .DIADI(B_write_data_low),                 // 16-bit input: A port data/LSB data
      .DIPADIP(),             // 2-bit input: A port parity/LSB parity
      // Port B Address/Control Signals: 14-bit (each) input: Port B address and control signals (write port
      // when RAM_MODE="SDP")
      .ADDRBWRADDR(write_address),     // 14-bit input: B port address/Write address
      .CLKBWRCLK(clk),         // 1-bit input: B port clock/Write clock
      .ENBWREN(1'b1),             // 1-bit input: B port enable/Write enable
      .REGCEB(),               // 1-bit input: B port register enable
      .RSTRAMB(),             // 1-bit input: B port set/reset
      .RSTREGB(),             // 1-bit input: B port register set/reset
      .WEBWE(write_enable),                 // 4-bit input: B port write enable/Write enable
      // Port B Data: 16-bit (each) input: Port B data
      .DIBDI(B_write_data_upper),                 // 16-bit input: B port data/MSB data
      .DIPBDIP()              // 2-bit input: B port parity/MSB parity
   );

   // End of RAMB18E1_inst instantiation

    endmodule
					
					
				
				